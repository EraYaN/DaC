configuration draw_rect_synthesised_cfg of draw_rect is
   for synthesised
   end for;
end draw_rect_synthesised_cfg;


