configuration rambank_synthesised_cfg of rambank is
   for synthesised
      for all: ramword use configuration work.ramword_behaviour_cfg;
      end for;
   end for;
end rambank_synthesised_cfg;


