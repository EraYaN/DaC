library IEEE;
use IEEE.std_logic_1164.ALL;
use work.parameter_def.ALL;

architecture behaviour of set_pixel is

begin
if(enable = '0')
color <= 'Z';
x0 <= 'Z';
y0 <= 'Z';
x1 <= 'Z';
y1 <= 'Z';
end if
if(enable = '1')



end process;

end behaviour;




