configuration rambank_behaviour_cfg of rambank is
   for behaviour
      for all: ramword use configuration work.ramword_behaviour_cfg;
      end for;
   end for;
end rambank_behaviour_cfg;


