configuration pwm_gen_behaviour_cfg of pwm_gen is
   for behaviour
   end for;
end pwm_gen_behaviour_cfg;


