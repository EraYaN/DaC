configuration draw_pixel_extracted_cfg of draw_pixel is
   for extracted
   end for;
end draw_pixel_extracted_cfg;


