library IEEE;
use IEEE.std_logic_1164.ALL;

PACKAGE ram_params IS
constant N : INTEGER;
END ram_params;

PACKAGE BODY ram_params IS
constant N : INTEGER:=16;
END ram_params;


