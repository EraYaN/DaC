library IEEE;
use IEEE.std_logic_1164.ALL;
use work.parameter_def.ALL;

entity decoder is
	port (
		--Clock/reset
		clk		: in	std_logic;						--Clock
		rst		: in	std_logic;						--Reset
		--SPI-interface interaction
		di		: in	std_logic_vector(7 downto 0);	--Data In
		do		: out	std_logic_vector(7 downto 0);	--Data Out
		dav		: in	std_logic;						--Data Available in SPI interface, commence data sampling
		rts		: out	std_logic;						--Ready To Send to SPI interface
		--Draw data
		x0		: out	std_logic_vector(7 downto 0);	--Entity x0 coord
		x1		: out	std_logic_vector(7 downto 0);	--Entity x1 coord
		y0		: out	std_logic_vector(7 downto 0);	--Entity y0 coord
		y1		: out	std_logic_vector(7 downto 0);	--Entity y1 coord
		col		: out	std_logic_vector(3 downto 0);	--Entity Color
		dwr		: in	std_logic;						--Draw Ready
		en		: out	std_logic_vector((NumDrawModules - 1) downto 0); --Draw Module Enabled
		--Internal registers
		id		: out	std_logic;						--Register id/address
		val		: out	std_logic;						--Value
		set		: out	std_logic						--Set
	);
end entity decoder;