library IEEE;
use IEEE.std_logic_1164.ALL;

entity vgacontrol_tb is
end vgacontrol_tb;


