configuration ramcontroller_behaviour_cfg of ramcontroller is
   for behaviour
   end for;
end ramcontroller_behaviour_cfg;


