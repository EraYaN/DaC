configuration alu_extracted_cfg of alu is
   for extracted
   end for;
end alu_extracted_cfg;


