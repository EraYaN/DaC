configuration alu_synthesised_cfg of alu is
   for synthesised
   end for;
end alu_synthesised_cfg;


