configuration alu_behaviour_cfg of alu is
   for behaviour
   end for;
end alu_behaviour_cfg;


