library IEEE;
use IEEE.std_logic_1164.ALL;
use ieee.numeric_std.all;


entity tb is
end tb;


