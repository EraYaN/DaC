configuration draw_pixel_behaviour_cfg of draw_pixel is
   for behaviour
   end for;
end draw_pixel_behaviour_cfg;


