configuration ramword_tb_behaviour_cfg of ramword_tb is
   for behaviour
      for all: ramword use configuration work.ramword_behaviour_cfg;
      end for;
   end for;
end ramword_tb_behaviour_cfg;


