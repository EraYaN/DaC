configuration draw_pixel_synthesised_cfg of draw_pixel is
   for synthesised
   end for;
end draw_pixel_synthesised_cfg;


