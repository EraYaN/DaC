configuration draw_rect_tb_behaviour_cfg of draw_rect_tb is
   for behaviour
      for all: draw_rect use configuration work.draw_rect_behaviour_cfg;
      end for;
   end for;
end draw_rect_tb_behaviour_cfg;


