library IEEE;
use IEEE.std_logic_1164.ALL;

entity draw_rect_tb is
end draw_rect_tb;