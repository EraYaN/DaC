library IEEE;
use IEEE.std_logic_1164.ALL;

entity draw_line_tb is
end draw_line_tb;