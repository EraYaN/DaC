configuration vgacontroller_behaviour_cfg of vgacontroller is
   for behaviour
   end for;
end vgacontroller_behaviour_cfg;


