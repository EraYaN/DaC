configuration rammux_synthesised_cfg of rammux is
   for synthesised
   end for;
end rammux_synthesised_cfg;


