library IEEE;
use IEEE.std_logic_1164.ALL;

entity decoder_tb is
end decoder_tb;