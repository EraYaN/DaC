* H:\GitHub\DaC\docs\opdracht 4\unified-model-parameters\NMOS.sch

* Schematics Version 9.1 - Web Update 1
* Mon Sep 30 10:45:51 2013



** Analysis setup **
.DC LIN V_V1 0 7 0.05 
.STEP LIN V_V2 0 5 1 
.OP 
.LIB "h:\Desktop\ModelLibEPO3.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "NMOS.net"
.INC "NMOS.als"


.probe


.END
