library IEEE;
use IEEE.std_logic_1164.ALL;

entity draw_pixel_tb is
end draw_pixel_tb;


