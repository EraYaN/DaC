library IEEE;
use IEEE.std_logic_1164.ALL;

entity rambank_tb is
end rambank_tb;


