configuration rammux_behaviour_cfg of rammux is
   for behaviour
   end for;
end rammux_behaviour_cfg;


