library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.ALL;

library work;
PACKAGE ramlib IS
constant WORDS : INTEGER:=8; -- number of words
constant ADRESSLINES: INTEGER:=3; -- numer of adresslines
constant WORDSIZE : INTEGER:=8; -- word size
END ramlib;

PACKAGE BODY ramlib IS


END ramlib;
















































