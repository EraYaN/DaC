library IEEE;
use IEEE.std_logic_1164.ALL;

entity ramword_tb is
end ramword_tb;


