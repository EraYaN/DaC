configuration pwm_gen_synthesised_cfg of pwm_gen is
   for synthesised
   end for;
end pwm_gen_synthesised_cfg;


