configuration draw_rect_behaviour_cfg of draw_rect is
   for behaviour
   end for;
end draw_rect_behaviour_cfg;


