configuration ramword_behaviour_cfg of ramword is
   for behaviour
   end for;
end ramword_behaviour_cfg;


