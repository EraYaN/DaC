library IEEE;
use IEEE.std_logic_1164.ALL;

PACKAGE parameter_def IS
	constant NumDrawModules : INTEGER;
	constant SizeX : INTEGER;
	constant SizeY : INTEGER;
	constant SizeMaxStageReg : INTEGER;
	constant NumStateReg : INTEGER;
	constant SizeRAMData : INTEGER;
	constant SizeRAMAddr : INTEGER;
	constant SizeColor : INTEGER;
END parameter_def;

PACKAGE BODY parameter_def IS
	constant NumDrawModules : INTEGER := 4; -- 0: pixel; 1: square; 2: line; 3: circle;
	constant SizeX : INTEGER := 8;
	constant SizeY : INTEGER := 7;
	constant SizeMaxStageReg : INTEGER := 1;
	constant NumStateReg : INTEGER := 1;
	constant SizeRAMData : INTEGER := 4;
	constant SizeRAMAddr : INTEGER := 16;
	constant SizeColor : INTEGER := 4;
END parameter_def;