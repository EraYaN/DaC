configuration spi_logic_cfg of spi is
   for logic
   end for;
end spi_logic_cfg;


