library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.ALL;

library work;
PACKAGE ramlib IS
constant WORDS : INTEGER:=4; -- number of words
constant ADRESSLINES: INTEGER:=2; -- numer of adresslines
constant WORDSIZE : INTEGER:=4; -- word size
END ramlib;

PACKAGE BODY ramlib IS


END ramlib;

































