* H:\GitHub\DaC\docs\opdracht 4\unified-model-parameters\resource\NMOS.sch

* Schematics Version 9.1 - Web Update 1
* Mon Oct 07 10:28:32 2013



** Analysis setup **
.DC LIN V_V1 0 7 0.05 
.STEP LIN V_V2 1 5 0.2 
.LIB "h:\Desktop\ModelLibEPO3.lib"
.LIB "h:\Desktop\ModelLibEPO3.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "NMOS.net"
.INC "NMOS.als"


.probe


.END
