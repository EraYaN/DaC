configuration ramcontroller_synthesised_cfg of ramcontroller is
   for synthesised
   end for;
end ramcontroller_synthesised_cfg;


